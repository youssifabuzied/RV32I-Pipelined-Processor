module InstMem (input [5:0] addr, output [31:0] data_out);
 reg [31:0] mem [0:63];
initial begin
mem[0]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0//added to be skipped since PC starts with 4 after reset 
mem[1]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0) 
mem[2]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[3]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[4]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[5]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0) 
mem[6]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[7]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[8]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[9]=32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0) 
mem[10]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[11]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[12]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[13]=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2 
mem[14]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[15]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[16]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[17]=32'b0_000001_00011_00100_000_0000_0_1100011; //beq x4, x3, 16
mem[18]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[19]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[20]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[21]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2 
mem[22]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[23]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[24]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[25]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2 
mem[26]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[27]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[28]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
mem[29]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0) 
mem[30]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[31]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[32]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[33]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
mem[34]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[35]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[36]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[37]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1 
mem[38]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[39]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[40]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[41]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2 
mem[42]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[43]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[44]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[45]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2 
mem[46]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[47]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[48]=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
mem[49]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
//mem[0] = 32'h028880B7;
//mem[1] = 32'h02888117;
//mem[2] = 32'h002081B3;
//mem[3] = 32'h00508213;
//mem[4] = 32'h0A020463;
//mem[5] = 32'h00400A6F;
//mem[6] = 32'h08119C63;
//mem[7] = 32'h00400A6F;
//mem[8] = 32'h0841C863;
//mem[9] = 32'h00400A6F;
//mem[10] = 32'h0811D463;
//mem[11] = 32'h0811E663;
//mem[12] = 32'h00400A6F;
//mem[13] = 32'h00000013;
//mem[14] = 32'h0011F463;
//mem[15] = 32'h00000013;
//mem[16] = 32'h00100283;
//mem[17] = 32'h00601303;
//mem[18] = 32'h00802383;
//mem[19] = 32'h00104403;
//mem[20] = 32'h00605483;
//mem[21] = 32'h00500723;
//mem[22] = 32'h00601923;
//mem[23] = 32'h00702A23;
//mem[24] = 32'h0010A593;
//mem[25] = 32'h0010B613;
//mem[26] = 32'h0010C693;
//mem[27] = 32'h0010E713;
//mem[28] = 32'h0010F793;
//mem[29] = 32'h00109813;
//mem[30] = 32'h0010D893;
//mem[31] = 32'h4010D913;
//mem[32] = 32'h00208533;
//mem[33] = 32'h402085B3;
//mem[34] = 32'h00209633;
//mem[35] = 32'h0020A6B3;
//mem[36] = 32'h0020B733;
//mem[37] = 32'h0020C7B3;
//mem[38] = 32'h0020D833;
//mem[39] = 32'h4020D8B3;
//mem[40] = 32'h0020E933;
//mem[41] = 32'h0020F4B3;
//mem[42] = 32'h0000000F;
//mem[43] = 32'h00000073;
//mem[44] = 32'h002181B3;
//mem[45] = 32'h004A0067;
//mem[46] = 32'h02302023;
//mem[47] = 32'h00100073;
//        mem[0]=32'h0x00508093;  // addi x1, x1, 5
//        mem[1]=32'h0x00108463;  // addi x2, x2, -4
//        mem[2]=32'h0x00510113;  // beq x1, x1, 8
//        mem[3]=32'h0x00218193;  // addi x3, x0, 10
//        mem[4]=32'h00b00213;  //  addi x4 x0 11
//        mem[5]=32'h00209463;  //  bne x1 x2    
//        mem[6]=32'h00a00193;  //  addi x3 x0 10
//        mem[7]=32'h00c00213;  //  addi x4 x0 12
//        mem[8]=32'h0020d463;  //  bge x1 x2 8  
//        mem[9]=32'h00a00193;  //  addi x3 x0 10
//       mem[10]=32'h00d00213; //  addi x4 x0 13
//       mem[11]=32'h0020e463; //  bltu x1 x2 8
//       mem[12]=32'h00a00193; //  addi x3 x0 10
//       mem[13]=32'h00e00213; //  addi x4 x0 14
//       mem[14]=32'h00114463; //  blt x2, x1, 8
//       mem[15]=32'h00a00193; //  addi x3, x0, 10
//       mem[16]=32'h00f00213; //  addi x4, x0, 15
//       mem[17]=32'h00117463; //  bgeu x2, x1, 8
//       mem[18]=32'h00a00193; //  addi x3, x0, 10
//       mem[19]=32'h01000213; //  addi x4, x0, 16
// mem[0]=32'b11111111101000000000000010010011 ; //lw x1, 0(x0)
 //mem[1]=32'b11111111101100000000000100010011 ; //lw x2, 4(x0)
// mem[2]=32'b00000000000100010010000110110011 ; //lw x3, 8(x0)
 //mem[3]=32'b00000110010000011000000101100111 ; //or x4, x1, x2

// mem[4]=32'b00000000000100011000000110010011; //beq x4, x3, 4
 
// mem[5]=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
// mem[6]=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
// mem[7]=32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
// mem[8]=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
// mem[9]=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
// mem[10]=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
// mem[11]=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
// mem[12]=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1*/
 

//        mem[0] = 32'b00000000000000000010001010000011; // lw lw x5, 0(x0)
//        mem[1] = 32'b00000000000000000001001100000011; //lh x6, 0(x0)
//        mem[2] = 32'b00000000000000000101001110000011;//lhu x7, 0(x0)
//        mem[3] = 32'b00000000000000000000111000000011; // lb x28,0(x0) 
//        mem[4] = 32'b00000000000000000100111010000011; // lbu x29, 0(x0)
//        mem[5] = 32'b00000000011000000010010000100011; // sw x6, 8(x0)
//        mem[6] = 32'b00000000011000000001010100100011; // sh x6, 10(x0)
//        mem[7] = 32'b00000000011000000000100010100011; // sb x6, 17(x0)
//        mem[8] = 32'b00000000100000000010010010000011; // lw x9, 8(x0)
//        mem[9] = 32'b00000000110000000010100100000011; //lw x18, 12(x0)
//        mem[10] = 32'b00000001000000000010100110000011; // lw x19, 16(x0)

end 
 assign data_out = mem[addr];
endmodule
